module Adder_4bits (input [3:0] A,B, output [3:0] C);
assign C = A + B;
endmodule